`define DISPLAY 1
`define NUMTAGTABLES 4
`define TABLESIZE 1024
`define BIMODALSIZE 2048
`define TAG1_SIZE 8
`define TAG2_SIZE 9
`define GEOMETRIC1 5
`define GEOMETRIC2 15
`define GEOMETRIC3 44
`define GEOMETRIC4 130
`define BIMODAL_LEN 11
`define TABLE_LEN 10
`define PHR_LEN 32

`define traceSize 3771697
